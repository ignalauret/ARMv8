module signext
  (input logic [31:0] a,
   output logic [63:0] y);

  always_comb 
    begin
      casez (a[31:21])
        11'b111_1100_00?0: y = { {56{a[20]}}, a[19:12] };
        11'b101_1010_0???: y = { {45{a[23]}}, a[22:5]  };
        default: y = 64'h0000000000000000;
      endcase
    end

endmodule

/*

  #OPCODE = 11 bits

  +---------------+--------+-----------------------------+-------------+--------+
  |  INSTRUCTION  |  TYPE  |           OPCODE            |  INDMEDIATE |  SIGN  |
  +---------------+--------+-----------------------------+-------------+--------+
  |     LDUR      |   D    |  0x7C2,     b111_1100_0010  |   [20:12]   |   Yes  |
  +---------------+--------+-----------------------------+-------------+--------+
  |     STUR      |   D    |  0x7C0,     b111_1100_0000  |   [20:12]   |   Yes  |
  +---------------+--------+-----------------------------+-------------+--------+
  |     CBZ       |   CB   |  0x5A0-5A7, b101_1010_0XXX  |   [23:5]    |   Yes  |
  +---------------+--------+-----------------------------+-------------+--------+

*/
